module ALU (input alu_op,
            input alu_in_1,
            input alu_in_2,
            output reg alu_result,
            output reg alu_bcond);  

endmodule