module ImmediateGenerator (input part_of_inst,
                           output reg imm_gen_out);  

endmodule
