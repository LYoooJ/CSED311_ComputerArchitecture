module alu (input alu_op, 
            input alu_in_1,
            input alu_in_2,
            output alu_result,
            output alu_bcond);

endmodule