module ALUControlUnit (input part_of_inst,
                       output reg alu_op);  
  
endmodule
