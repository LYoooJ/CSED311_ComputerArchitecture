module pc(.reset(),clk(),next_pc());


endmodule