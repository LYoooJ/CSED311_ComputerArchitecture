module alu () ();

endmodule