module alu_control_unit(part_of_inst(),alu_op());



endmodule
